LIBRARY library IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY Vending_Machine IS
    PORT ();
END Vending_Machine;

ARCHITECTURE Behavioral OF Vending_Machine IS

BEGIN

END Behavioral;